diffBuf_inst : diffBuf PORT MAP (
		datain	 => datain_sig,
		dataout	 => dataout_sig,
		dataout_b	 => dataout_b_sig
	);
